-- Synthesis only
library ieee;
use ieee.std_logic_1164.all;
use ieee.fixed_pkg.all; 

use work.rnn_pkg.all;

entity tanh_lut is
    port (
        x : in acc_t;
        y : out tanh_t
    );
end entity tanh_lut;

architecture behav of tanh_lut is
begin    
    process (x) is
        variable x_addr : std_logic_vector(7 downto 0);
        variable y_ram : tanh_t;
    begin
        x_addr := to_slv(x(1 downto -6));

        case x_addr is
            when "00000000" => y_ram := to_sfixed(0.0, y'high, y'low);
            when "00000001" => y_ram := to_sfixed(0.01556396484375, y'high, y'low);
            when "00000010" => y_ram := to_sfixed(0.03118896484375, y'high, y'low);
            when "00000011" => y_ram := to_sfixed(0.04681396484375, y'high, y'low);
            when "00000100" => y_ram := to_sfixed(0.0623779296875, y'high, y'low);
            when "00000101" => y_ram := to_sfixed(0.07794189453125, y'high, y'low);
            when "00000110" => y_ram := to_sfixed(0.09344482421875, y'high, y'low);
            when "00000111" => y_ram := to_sfixed(0.10888671875, y'high, y'low);
            when "00001000" => y_ram := to_sfixed(0.12432861328125, y'high, y'low);
            when "00001001" => y_ram := to_sfixed(0.1396484375, y'high, y'low);
            when "00001010" => y_ram := to_sfixed(0.15496826171875, y'high, y'low);
            when "00001011" => y_ram := to_sfixed(0.170166015625, y'high, y'low);
            when "00001100" => y_ram := to_sfixed(0.185302734375, y'high, y'low);
            when "00001101" => y_ram := to_sfixed(0.2003173828125, y'high, y'low);
            when "00001110" => y_ram := to_sfixed(0.21527099609375, y'high, y'low);
            when "00001111" => y_ram := to_sfixed(0.23016357421875, y'high, y'low);
            when "00010000" => y_ram := to_sfixed(0.244873046875, y'high, y'low);
            when "00010001" => y_ram := to_sfixed(0.259521484375, y'high, y'low);
            when "00010010" => y_ram := to_sfixed(0.2740478515625, y'high, y'low);
            when "00010011" => y_ram := to_sfixed(0.28839111328125, y'high, y'low);
            when "00010100" => y_ram := to_sfixed(0.30267333984375, y'high, y'low);
            when "00010101" => y_ram := to_sfixed(0.31683349609375, y'high, y'low);
            when "00010110" => y_ram := to_sfixed(0.330810546875, y'high, y'low);
            when "00010111" => y_ram := to_sfixed(0.3446044921875, y'high, y'low);
            when "00011000" => y_ram := to_sfixed(0.35833740234375, y'high, y'low);
            when "00011001" => y_ram := to_sfixed(0.37188720703125, y'high, y'low);
            when "00011010" => y_ram := to_sfixed(0.38525390625, y'high, y'low);
            when "00011011" => y_ram := to_sfixed(0.39849853515625, y'high, y'low);
            when "00011100" => y_ram := to_sfixed(0.41156005859375, y'high, y'low);
            when "00011101" => y_ram := to_sfixed(0.4244384765625, y'high, y'low);
            when "00011110" => y_ram := to_sfixed(0.4371337890625, y'high, y'low);
            when "00011111" => y_ram := to_sfixed(0.44970703125, y'high, y'low);
            when "00100000" => y_ram := to_sfixed(0.46209716796875, y'high, y'low);
            when "00100001" => y_ram := to_sfixed(0.47430419921875, y'high, y'low);
            when "00100010" => y_ram := to_sfixed(0.486328125, y'high, y'low);
            when "00100011" => y_ram := to_sfixed(0.4981689453125, y'high, y'low);
            when "00100100" => y_ram := to_sfixed(0.50982666015625, y'high, y'low);
            when "00100101" => y_ram := to_sfixed(0.52130126953125, y'high, y'low);
            when "00100110" => y_ram := to_sfixed(0.53253173828125, y'high, y'low);
            when "00100111" => y_ram := to_sfixed(0.54364013671875, y'high, y'low);
            when "00101000" => y_ram := to_sfixed(0.5545654296875, y'high, y'low);
            when "00101001" => y_ram := to_sfixed(0.5653076171875, y'high, y'low);
            when "00101010" => y_ram := to_sfixed(0.5758056640625, y'high, y'low);
            when "00101011" => y_ram := to_sfixed(0.586181640625, y'high, y'low);
            when "00101100" => y_ram := to_sfixed(0.5963134765625, y'high, y'low);
            when "00101101" => y_ram := to_sfixed(0.6063232421875, y'high, y'low);
            when "00101110" => y_ram := to_sfixed(0.6160888671875, y'high, y'low);
            when "00101111" => y_ram := to_sfixed(0.625732421875, y'high, y'low);
            when "00110000" => y_ram := to_sfixed(0.6351318359375, y'high, y'low);
            when "00110001" => y_ram := to_sfixed(0.64434814453125, y'high, y'low);
            when "00110010" => y_ram := to_sfixed(0.65338134765625, y'high, y'low);
            when "00110011" => y_ram := to_sfixed(0.6622314453125, y'high, y'low);
            when "00110100" => y_ram := to_sfixed(0.67095947265625, y'high, y'low);
            when "00110101" => y_ram := to_sfixed(0.679443359375, y'high, y'low);
            when "00110110" => y_ram := to_sfixed(0.687744140625, y'high, y'low);
            when "00110111" => y_ram := to_sfixed(0.6959228515625, y'high, y'low);
            when "00111000" => y_ram := to_sfixed(0.703857421875, y'high, y'low);
            when "00111001" => y_ram := to_sfixed(0.711669921875, y'high, y'low);
            when "00111010" => y_ram := to_sfixed(0.71929931640625, y'high, y'low);
            when "00111011" => y_ram := to_sfixed(0.72674560546875, y'high, y'low);
            when "00111100" => y_ram := to_sfixed(0.73406982421875, y'high, y'low);
            when "00111101" => y_ram := to_sfixed(0.74114990234375, y'high, y'low);
            when "00111110" => y_ram := to_sfixed(0.74810791015625, y'high, y'low);
            when "00111111" => y_ram := to_sfixed(0.75494384765625, y'high, y'low);
            when "01000000" => y_ram := to_sfixed(0.76153564453125, y'high, y'low);
            when "01000001" => y_ram := to_sfixed(0.76806640625, y'high, y'low);
            when "01000010" => y_ram := to_sfixed(0.77435302734375, y'high, y'low);
            when "01000011" => y_ram := to_sfixed(0.78057861328125, y'high, y'low);
            when "01000100" => y_ram := to_sfixed(0.78656005859375, y'high, y'low);
            when "01000101" => y_ram := to_sfixed(0.79248046875, y'high, y'low);
            when "01000110" => y_ram := to_sfixed(0.7982177734375, y'high, y'low);
            when "01000111" => y_ram := to_sfixed(0.8038330078125, y'high, y'low);
            when "01001000" => y_ram := to_sfixed(0.80926513671875, y'high, y'low);
            when "01001001" => y_ram := to_sfixed(0.8145751953125, y'high, y'low);
            when "01001010" => y_ram := to_sfixed(0.81976318359375, y'high, y'low);
            when "01001011" => y_ram := to_sfixed(0.8248291015625, y'high, y'low);
            when "01001100" => y_ram := to_sfixed(0.82977294921875, y'high, y'low);
            when "01001101" => y_ram := to_sfixed(0.8345947265625, y'high, y'low);
            when "01001110" => y_ram := to_sfixed(0.8392333984375, y'high, y'low);
            when "01001111" => y_ram := to_sfixed(0.84381103515625, y'high, y'low);
            when "01010000" => y_ram := to_sfixed(0.8482666015625, y'high, y'low);
            when "01010001" => y_ram := to_sfixed(0.85260009765625, y'high, y'low);
            when "01010010" => y_ram := to_sfixed(0.8568115234375, y'high, y'low);
            when "01010011" => y_ram := to_sfixed(0.86090087890625, y'high, y'low);
            when "01010100" => y_ram := to_sfixed(0.8648681640625, y'high, y'low);
            when "01010101" => y_ram := to_sfixed(0.8687744140625, y'high, y'low);
            when "01010110" => y_ram := to_sfixed(0.87255859375, y'high, y'low);
            when "01010111" => y_ram := to_sfixed(0.876220703125, y'high, y'low);
            when "01011000" => y_ram := to_sfixed(0.87982177734375, y'high, y'low);
            when "01011001" => y_ram := to_sfixed(0.88330078125, y'high, y'low);
            when "01011010" => y_ram := to_sfixed(0.88665771484375, y'high, y'low);
            when "01011011" => y_ram := to_sfixed(0.88995361328125, y'high, y'low);
            when "01011100" => y_ram := to_sfixed(0.8931884765625, y'high, y'low);
            when "01011101" => y_ram := to_sfixed(0.89630126953125, y'high, y'low);
            when "01011110" => y_ram := to_sfixed(0.8992919921875, y'high, y'low);
            when "01011111" => y_ram := to_sfixed(0.90228271484375, y'high, y'low);
            when "01100000" => y_ram := to_sfixed(0.90509033203125, y'high, y'low);
            when "01100001" => y_ram := to_sfixed(0.90789794921875, y'high, y'low);
            when "01100010" => y_ram := to_sfixed(0.91058349609375, y'high, y'low);
            when "01100011" => y_ram := to_sfixed(0.9132080078125, y'high, y'low);
            when "01100100" => y_ram := to_sfixed(0.915771484375, y'high, y'low);
            when "01100101" => y_ram := to_sfixed(0.91827392578125, y'high, y'low);
            when "01100110" => y_ram := to_sfixed(0.92071533203125, y'high, y'low);
            when "01100111" => y_ram := to_sfixed(0.92303466796875, y'high, y'low);
            when "01101000" => y_ram := to_sfixed(0.92529296875, y'high, y'low);
            when "01101001" => y_ram := to_sfixed(0.92755126953125, y'high, y'low);
            when "01101010" => y_ram := to_sfixed(0.9296875, y'high, y'low);
            when "01101011" => y_ram := to_sfixed(0.9317626953125, y'high, y'low);
            when "01101100" => y_ram := to_sfixed(0.93377685546875, y'high, y'low);
            when "01101101" => y_ram := to_sfixed(0.935791015625, y'high, y'low);
            when "01101110" => y_ram := to_sfixed(0.93768310546875, y'high, y'low);
            when "01101111" => y_ram := to_sfixed(0.93951416015625, y'high, y'low);
            when "01110000" => y_ram := to_sfixed(0.94134521484375, y'high, y'low);
            when "01110001" => y_ram := to_sfixed(0.943115234375, y'high, y'low);
            when "01110010" => y_ram := to_sfixed(0.94482421875, y'high, y'low);
            when "01110011" => y_ram := to_sfixed(0.94647216796875, y'high, y'low);
            when "01110100" => y_ram := to_sfixed(0.94805908203125, y'high, y'low);
            when "01110101" => y_ram := to_sfixed(0.9495849609375, y'high, y'low);
            when "01110110" => y_ram := to_sfixed(0.95111083984375, y'high, y'low);
            when "01110111" => y_ram := to_sfixed(0.95257568359375, y'high, y'low);
            when "01111000" => y_ram := to_sfixed(0.95404052734375, y'high, y'low);
            when "01111001" => y_ram := to_sfixed(0.95538330078125, y'high, y'low);
            when "01111010" => y_ram := to_sfixed(0.95672607421875, y'high, y'low);
            when "01111011" => y_ram := to_sfixed(0.95806884765625, y'high, y'low);
            when "01111100" => y_ram := to_sfixed(0.95928955078125, y'high, y'low);
            when "01111101" => y_ram := to_sfixed(0.96051025390625, y'high, y'low);
            when "01111110" => y_ram := to_sfixed(0.96173095703125, y'high, y'low);
            when "01111111" => y_ram := to_sfixed(0.962890625, y'high, y'low);
            when "10000000" => y_ram := to_sfixed(0.9639892578125, y'high, y'low);
            when "10000001" => y_ram := to_sfixed(0.965087890625, y'high, y'low);
            when "10000010" => y_ram := to_sfixed(0.96612548828125, y'high, y'low);
            when "10000011" => y_ram := to_sfixed(0.9671630859375, y'high, y'low);
            when "10000100" => y_ram := to_sfixed(0.9681396484375, y'high, y'low);
            when "10000101" => y_ram := to_sfixed(0.9691162109375, y'high, y'low);
            when "10000110" => y_ram := to_sfixed(0.97003173828125, y'high, y'low);
            when "10000111" => y_ram := to_sfixed(0.970947265625, y'high, y'low);
            when "10001000" => y_ram := to_sfixed(0.97186279296875, y'high, y'low);
            when "10001001" => y_ram := to_sfixed(0.97271728515625, y'high, y'low);
            when "10001010" => y_ram := to_sfixed(0.9735107421875, y'high, y'low);
            when "10001011" => y_ram := to_sfixed(0.97430419921875, y'high, y'low);
            when "10001100" => y_ram := to_sfixed(0.97509765625, y'high, y'low);
            when "10001101" => y_ram := to_sfixed(0.97589111328125, y'high, y'low);
            when "10001110" => y_ram := to_sfixed(0.97662353515625, y'high, y'low);
            when "10001111" => y_ram := to_sfixed(0.977294921875, y'high, y'low);
            when "10010000" => y_ram := to_sfixed(0.97796630859375, y'high, y'low);
            when "10010001" => y_ram := to_sfixed(0.9786376953125, y'high, y'low);
            when "10010010" => y_ram := to_sfixed(0.97930908203125, y'high, y'low);
            when "10010011" => y_ram := to_sfixed(0.97991943359375, y'high, y'low);
            when "10010100" => y_ram := to_sfixed(0.98052978515625, y'high, y'low);
            when "10010101" => y_ram := to_sfixed(0.98114013671875, y'high, y'low);
            when "10010110" => y_ram := to_sfixed(0.981689453125, y'high, y'low);
            when "10010111" => y_ram := to_sfixed(0.9822998046875, y'high, y'low);
            when "10011000" => y_ram := to_sfixed(0.9827880859375, y'high, y'low);
            when "10011001" => y_ram := to_sfixed(0.98333740234375, y'high, y'low);
            when "10011010" => y_ram := to_sfixed(0.98382568359375, y'high, y'low);
            when "10011011" => y_ram := to_sfixed(0.98431396484375, y'high, y'low);
            when "10011100" => y_ram := to_sfixed(0.98480224609375, y'high, y'low);
            when "10011101" => y_ram := to_sfixed(0.98529052734375, y'high, y'low);
            when "10011110" => y_ram := to_sfixed(0.9857177734375, y'high, y'low);
            when "10011111" => y_ram := to_sfixed(0.98614501953125, y'high, y'low);
            when "10100000" => y_ram := to_sfixed(0.986572265625, y'high, y'low);
            when "10100001" => y_ram := to_sfixed(0.98699951171875, y'high, y'low);
            when "10100010" => y_ram := to_sfixed(0.98736572265625, y'high, y'low);
            when "10100011" => y_ram := to_sfixed(0.98779296875, y'high, y'low);
            when "10100100" => y_ram := to_sfixed(0.9881591796875, y'high, y'low);
            when "10100101" => y_ram := to_sfixed(0.988525390625, y'high, y'low);
            when "10100110" => y_ram := to_sfixed(0.98883056640625, y'high, y'low);
            when "10100111" => y_ram := to_sfixed(0.98919677734375, y'high, y'low);
            when "10101000" => y_ram := to_sfixed(0.989501953125, y'high, y'low);
            when "10101001" => y_ram := to_sfixed(0.9898681640625, y'high, y'low);
            when "10101010" => y_ram := to_sfixed(0.99017333984375, y'high, y'low);
            when "10101011" => y_ram := to_sfixed(0.990478515625, y'high, y'low);
            when "10101100" => y_ram := to_sfixed(0.99072265625, y'high, y'low);
            when "10101101" => y_ram := to_sfixed(0.99102783203125, y'high, y'low);
            when "10101110" => y_ram := to_sfixed(0.9913330078125, y'high, y'low);
            when "10101111" => y_ram := to_sfixed(0.9915771484375, y'high, y'low);
            when "10110000" => y_ram := to_sfixed(0.9918212890625, y'high, y'low);
            when "10110001" => y_ram := to_sfixed(0.9920654296875, y'high, y'low);
            when "10110010" => y_ram := to_sfixed(0.9923095703125, y'high, y'low);
            when "10110011" => y_ram := to_sfixed(0.9925537109375, y'high, y'low);
            when "10110100" => y_ram := to_sfixed(0.9927978515625, y'high, y'low);
            when "10110101" => y_ram := to_sfixed(0.99298095703125, y'high, y'low);
            when "10110110" => y_ram := to_sfixed(0.99322509765625, y'high, y'low);
            when "10110111" => y_ram := to_sfixed(0.993408203125, y'high, y'low);
            when "10111000" => y_ram := to_sfixed(0.99365234375, y'high, y'low);
            when "10111001" => y_ram := to_sfixed(0.99383544921875, y'high, y'low);
            when "10111010" => y_ram := to_sfixed(0.9940185546875, y'high, y'low);
            when "10111011" => y_ram := to_sfixed(0.99420166015625, y'high, y'low);
            when "10111100" => y_ram := to_sfixed(0.994384765625, y'high, y'low);
            when "10111101" => y_ram := to_sfixed(0.99456787109375, y'high, y'low);
            when "10111110" => y_ram := to_sfixed(0.99468994140625, y'high, y'low);
            when "10111111" => y_ram := to_sfixed(0.994873046875, y'high, y'low);
            when "11000000" => y_ram := to_sfixed(0.9949951171875, y'high, y'low);
            when "11000001" => y_ram := to_sfixed(0.99517822265625, y'high, y'low);
            when "11000010" => y_ram := to_sfixed(0.99530029296875, y'high, y'low);
            when "11000011" => y_ram := to_sfixed(0.9954833984375, y'high, y'low);
            when "11000100" => y_ram := to_sfixed(0.99560546875, y'high, y'low);
            when "11000101" => y_ram := to_sfixed(0.9957275390625, y'high, y'low);
            when "11000110" => y_ram := to_sfixed(0.995849609375, y'high, y'low);
            when "11000111" => y_ram := to_sfixed(0.9959716796875, y'high, y'low);
            when "11001000" => y_ram := to_sfixed(0.99609375, y'high, y'low);
            when "11001001" => y_ram := to_sfixed(0.9962158203125, y'high, y'low);
            when "11001010" => y_ram := to_sfixed(0.996337890625, y'high, y'low);
            when "11001011" => y_ram := to_sfixed(0.9964599609375, y'high, y'low);
            when "11001100" => y_ram := to_sfixed(0.99658203125, y'high, y'low);
            when "11001101" => y_ram := to_sfixed(0.99664306640625, y'high, y'low);
            when "11001110" => y_ram := to_sfixed(0.99676513671875, y'high, y'low);
            when "11001111" => y_ram := to_sfixed(0.99688720703125, y'high, y'low);
            when "11010000" => y_ram := to_sfixed(0.9969482421875, y'high, y'low);
            when "11010001" => y_ram := to_sfixed(0.9970703125, y'high, y'low);
            when "11010010" => y_ram := to_sfixed(0.99713134765625, y'high, y'low);
            when "11010011" => y_ram := to_sfixed(0.99725341796875, y'high, y'low);
            when "11010100" => y_ram := to_sfixed(0.997314453125, y'high, y'low);
            when "11010101" => y_ram := to_sfixed(0.99737548828125, y'high, y'low);
            when "11010110" => y_ram := to_sfixed(0.99749755859375, y'high, y'low);
            when "11010111" => y_ram := to_sfixed(0.99755859375, y'high, y'low);
            when "11011000" => y_ram := to_sfixed(0.99761962890625, y'high, y'low);
            when "11011001" => y_ram := to_sfixed(0.9976806640625, y'high, y'low);
            when "11011010" => y_ram := to_sfixed(0.99774169921875, y'high, y'low);
            when "11011011" => y_ram := to_sfixed(0.99786376953125, y'high, y'low);
            when "11011100" => y_ram := to_sfixed(0.9979248046875, y'high, y'low);
            when "11011101" => y_ram := to_sfixed(0.99798583984375, y'high, y'low);
            when "11011110" => y_ram := to_sfixed(0.998046875, y'high, y'low);
            when "11011111" => y_ram := to_sfixed(0.99810791015625, y'high, y'low);
            when "11100000" => y_ram := to_sfixed(0.9981689453125, y'high, y'low);
            when "11100001" => y_ram := to_sfixed(0.99822998046875, y'high, y'low);
            when "11100010" => y_ram := to_sfixed(0.99822998046875, y'high, y'low);
            when "11100011" => y_ram := to_sfixed(0.998291015625, y'high, y'low);
            when "11100100" => y_ram := to_sfixed(0.99835205078125, y'high, y'low);
            when "11100101" => y_ram := to_sfixed(0.9984130859375, y'high, y'low);
            when "11100110" => y_ram := to_sfixed(0.99847412109375, y'high, y'low);
            when "11100111" => y_ram := to_sfixed(0.99853515625, y'high, y'low);
            when "11101000" => y_ram := to_sfixed(0.99853515625, y'high, y'low);
            when "11101001" => y_ram := to_sfixed(0.99859619140625, y'high, y'low);
            when "11101010" => y_ram := to_sfixed(0.9986572265625, y'high, y'low);
            when "11101011" => y_ram := to_sfixed(0.9986572265625, y'high, y'low);
            when "11101100" => y_ram := to_sfixed(0.99871826171875, y'high, y'low);
            when "11101101" => y_ram := to_sfixed(0.998779296875, y'high, y'low);
            when "11101110" => y_ram := to_sfixed(0.998779296875, y'high, y'low);
            when "11101111" => y_ram := to_sfixed(0.99884033203125, y'high, y'low);
            when "11110000" => y_ram := to_sfixed(0.99884033203125, y'high, y'low);
            when "11110001" => y_ram := to_sfixed(0.9989013671875, y'high, y'low);
            when "11110010" => y_ram := to_sfixed(0.9989013671875, y'high, y'low);
            when "11110011" => y_ram := to_sfixed(0.99896240234375, y'high, y'low);
            when "11110100" => y_ram := to_sfixed(0.9990234375, y'high, y'low);
            when "11110101" => y_ram := to_sfixed(0.9990234375, y'high, y'low);
            when "11110110" => y_ram := to_sfixed(0.9990234375, y'high, y'low);
            when "11110111" => y_ram := to_sfixed(0.99908447265625, y'high, y'low);
            when "11111000" => y_ram := to_sfixed(0.99908447265625, y'high, y'low);
            when "11111001" => y_ram := to_sfixed(0.9991455078125, y'high, y'low);
            when "11111010" => y_ram := to_sfixed(0.9991455078125, y'high, y'low);
            when "11111011" => y_ram := to_sfixed(0.99920654296875, y'high, y'low);
            when "11111100" => y_ram := to_sfixed(0.99920654296875, y'high, y'low);
            when "11111101" => y_ram := to_sfixed(0.99920654296875, y'high, y'low);
            when "11111110" => y_ram := to_sfixed(0.999267578125, y'high, y'low);
            when "11111111" => y_ram := to_sfixed(0.999267578125, y'high, y'low);
            when others => y_ram := to_sfixed(1.0, y'high, y'low);
        end case; 

        if x > 4.0 then
            y <= to_sfixed(1.0, y'high, y'low);
        elsif x >= 0.0 then
            y <= y_ram;
        elsif x >= -4.0 then
            y <= '1' & y_ram(0 downto y'low);
        else 
            y <= to_sfixed(-1.0, y'high, y'low);
        end if;
    end process;
        
                
end architecture behav;